class vec3fixed24x8;
    function new();
        
    endfunction //new()
endclass //vec3fixed24x8