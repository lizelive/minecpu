module mailbox_tb;
    mailbox #(int) mailbox = new(10);
endmodule